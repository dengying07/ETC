** Profile: "SCHEMATIC1-Bias"  [ C:\Users\deng\Desktop\ģ����\experiment\ʵ��4\bjt1-schematic1-bias.sim ] 

** Creating circuit file "bjt1-schematic1-bias.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of d:\orcad92\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 150ms 110ms 0.1m 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\BJT1-SCHEMATIC1.net" 


.END
