** Profile: "SCHEMATIC1-Bias"  [ D:\09300720075\d1101-schematic1-bias.sim ] 

** Creating circuit file "d1101-schematic1-bias.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1000u 0 1u 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\D1101-SCHEMATIC1.net" 


.END
