** Profile: "SCHEMATIC1-Bias"  [ C:\Users\deng\Desktop\ģ��\experiments\1_6_11_4jie-schematic1-bias.sim ] 

** Creating circuit file "1_6_11_4jie-schematic1-bias.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of d:\orcad92\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 100 1 100meg
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\1_6_11_4jie-SCHEMATIC1.net" 


.END
