LIBRARY ieee;
USE ieee.std_logic_1164.all;
Use IEEE.std_logic_unsigned.ALL;
ENTITY testbench IS
END ENTITY testbench;

ARCHITECTURE test OF testbench IS
	SIGNAL result_test: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL instuctionS_test: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL clk_test: STD_LOGIC;
	SIGNAL enable_test: STD_LOGIC;
BEGIN
	
g0:PROCESS	-- Define the clock
BEGIN
	clk_test<='1';
	WAIT FOR 25NS;
	clk_test<='0';
	WAIT FOR 25NS;
	END PROCESS;

g1:ENTITY work.microprocessor(behavior)
		PORT MAP (instructions=>instuctions_test,clk=>clk_test, enable=>enable_test,result=>result_test);
		instuctions_test <=B"00101100001000100000000000000000",		--r1+r2
			     B"00101100000001010000000000000000" AFTER 50NS,	--sum1+r5
			     B"00101100000001100000000000000000" AFTER 100NS,	--sum1+r6
			     B"00101100000010010000000000000000" AFTER 150NS,	--sum1+r9
			     B"00101100000010100000000000000000" AFTER 200NS,	--sum1+r10
			     B"00101100000011010000000000000000" AFTER 250NS,	--sum1+r13
			     B"00101100000011100000000000000000" AFTER 300NS,	--sum1+r14
			     B"00101100000100010000000000000000" AFTER 350NS,	--sum1+r17
			     B"00101100000100100000000000000000" AFTER 400NS,	--sum1+r18
			     B"00101100000101010000000000000000" AFTER 450NS,	--sum1+r21
			     B"00101100000100100000000000000000" AFTER 500NS,	--sum1+r22
			     B"00101100000110010000000000000000" AFTER 550NS,	--sum1+r25
			     B"00101100000110100000000000000000" AFTER 600NS,	--sum1+r26
			     B"00101100000111010000000000000000" AFTER 650NS,	--sum1+r29
			     B"00101100000111100000000000000000" AFTER 700NS,	--sum1+r30

			     B"00101100011001001111100000000000" AFTER 750NS,	--r3+r4
			     B"00101111111001111111100000000000" AFTER 800NS,	--sum2+r7
			     B"00101111111010001111100000000000" AFTER 850NS,	--sum2+r8
			     B"00101111111010111111100000000000" AFTER 900NS,	--sum2+r11
			     B"00101111111011001111100000000000" AFTER 950NS,	--sum2+r12
			     B"00101111111011111111100000000000" AFTER 1000NS,	--sum2+r15
			     B"00101111111100001111100000000000" AFTER 1050NS,	--sum2+r16
			     B"00101111111100111111100000000000" AFTER 1100NS,	--sum2+r19
			     B"00101111111101001111100000000000" AFTER 1150NS,	--sum2+r20
			     B"00101111111101111111100000000000" AFTER 1200NS,	--sum2+r23
			     B"00101111111110001111100000000000" AFTER 1250NS,	--sum2+r24
			     B"00101111111110111111100000000000" AFTER 1300NS,	--sum2+r27
			     B"00101111111111001111100000000000" AFTER 1350NS,	--sum2+r28

			     B"00011000000111111111100000000000" AFTER 1400NS;	--sum1-sum2
			
			     
				
				
	
END ARCHITECTURE test;