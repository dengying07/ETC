** Profile: "SCHEMATIC1-Bias"  [ C:\Users\deng\Desktop\ģ��\experiments\09300720075\1_6_5a-schematic1-bias.sim ] 

** Creating circuit file "1_6_5a-schematic1-bias.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of d:\orcad92\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN V_V3 -2 1.5 0.5 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\1_6_5a-SCHEMATIC1.net" 


.END
