** Profile: "SCHEMATIC1-Bias"  [ D:\09300720075\1_4_1-schematic1-bias.sim ] 

** Creating circuit file "1_4_1-schematic1-bias.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 5s 0 0.005 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\1_4_1-SCHEMATIC1.net" 


.END
