** Profile: "SCHEMATIC1-Bias"  [ D:\09300720075\1_3_1-schematic1-bias.sim ] 

** Creating circuit file "1_3_1-schematic1-bias.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 0.1m 0 0.0001m 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\1_3_1-SCHEMATIC1.net" 


.END
